// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 64-Bit Version 13.0 (Build Build 232 06/12/2013)
// Created on Tue Sep 10 02:55:15 2019
`timescale 1 ps / 1 ps

module LAB1_th;

	reg clk_sig;
	reg arstn_sig;
	reg we_sig;
	reg srstn_sig;
	reg [31:0] dat_sig;
	wire [31:0] dout_sig;

	LAB1 LAB1_inst
	(
		.we(we_sig),	// input  we_sig
		.srstn(srstn_sig),	// input  srstn_sig
		.clk(clk_sig),	// input  clk_sig
		.arstn(arstn_sig),	// input  arstn_sig
		.dat(dat_sig),	// input [31:0] dat_sig
		.dout(dout_sig) 	// output [31:0] dout_sig
	);

initial begin
	clk_sig =1'd1;
	forever #1 clk_sig = ~clk_sig;
end

initial begin
	arstn_sig =1'b1;
	we_sig =1'b1;
	
	#2 arstn_sig =1'b0;
	#2 arstn_sig =1'b1;
end

initial begin 
	srstn_sig =1'b1;
	
	#20 srstn_sig =1'b0;
	#5 srstn_sig =1'b1;
end

initial begin
	dat_sig = 32'h0;
	#10 dat_sig = 32'hdeadc0de;
	#30 dat_sig = 32'hdeadbeef;
end

initial begin
	#50 $stop();
end

endmodule	
	
