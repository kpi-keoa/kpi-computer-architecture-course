// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 32-bit Version 13.0 (Build Build 232 06/12/2013)
// Created on Sat Oct 12 17:48:46 20194

`timescale 1ns / 1ps

module alu_tb;

reg [31:0] i_a_sig;
reg [31:0] i_b_sig;
reg [1:0] i_alufunc_sig;
reg [2:0] i_opt_sig;

wire [31:0] o_result_sig;
wire o_zero_sig;
wire o_ovfl_sig;


alu alu_inst
(
	.i_a(i_a_sig),			// input [31:0] i_a_sig
	.i_b(i_b_sig),			// input [31:0] i_b_sig
	.i_opt(i_opt_sig),		// input [2:0] i_opt_sig
	.i_alufunc(i_alufunc_sig),	// input [1:0] i_alufunc_sig
	.o_result(o_result_sig),	// output [31:0] o_result_sig
	.o_zero(o_zero_sig),		// output  o_zero_sig
	.o_ovfl(o_ovfl_sig) 		// output  o_ovfl_sig
);

// Idea was taken from job of Kharchuk's Vadim

initial begin

	i_a_sig = 32'b00110011;		//add
	#20 i_a_sig = 32'b10101010; 	//mul
	#40 i_a_sig = 32'b11001010; 	//shif
	#50 i_a_sig = 32'b11100011; 	//logic	
	
end

initial begin

	i_b_sig = 32'b11001100;		//add
	#20 i_b_sig = 32'b00001111; 	//mul
	#40 i_b_sig = 32'b01010101;	//shift
	#50 i_b_sig = 32'b00101010; 	//logic

end


initial begin

	i_alufunc_sig = 2'b11;		// add
	#20 i_alufunc_sig = 2'b00;	// mul
	#40 i_alufunc_sig = 2'b10; 	// shift
	#50 i_alufunc_sig = 2'b01; 	// logic

end

initial begin
	i_opt_sig = 1'b0;		// test addsub
	#10 i_opt_sig = 1'b1;

	#10 i_opt_sig = 2'b00;		// Mult[63:32]
	#10 i_opt_sig = 2'b10;		// Mult[31:0]
	#10 i_opt_sig = 2'b01;		// Div
	#10 i_opt_sig = 2'b11;		// Module

	#10 i_opt_sig = 3'b000;		// Sll
	#10 i_opt_sig = 3'b001;		// SRl
	#10 i_opt_sig = 3'b010;		// ROL
	#10 i_opt_sig = 3'b011;		// ROR
	#10 i_opt_sig = 3'b111;		// SRA

	#10 i_opt_sig = 2'b01;	// &
	#10 i_opt_sig = 2'b10;	// |
	#10 i_opt_sig = 2'b00;	// ~( | )
	#10 i_opt_sig = 2'b11;	// ^
	
end

initial begin 
	#400 $stop();
end
endmodule


