// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 64-Bit Version 13.0 (Build Build 232 06/12/2013)
// Created on Tue Sep 24 21:21:42 2019

`timescale 1ns/1ps

module barrel_shifter_tb;

	reg  [2:0] bs_opsel_sig;
	reg  [4:0] shift_amount_sig;
	reg  [31:0] data_in_sig;
	wire [31:0] result_sig;

barrel_shifter barrel_shifter_inst
(
	.bs_opsel(bs_opsel_sig) ,	// input [2:0] bs_opsel_sig
	.shift_amount(shift_amount_sig) ,	// input [31:0] shift_amount_sig
	.data_in(data_in_sig) ,	// input [31:0] data_in_sig
	.result(result_sig) 	// output [31:0] result_sig
);

	initial begin 
		data_in_sig= 32'habcd1234;
		shift_amount_sig = 5'h4;
		
		bs_opsel_sig = 3'b000;		//shift left logical
		#10 bs_opsel_sig = 3'b001;	//rotate left
		#10 bs_opsel_sig = 3'b010;	//shift right logical
		#10 bs_opsel_sig = 3'b011;	//rotate right
		#10 bs_opsel_sig = 3'b111;	//shift right arithmetical]

		end

	initial begin
		#50 $stop();
		end


endmodule

