`define bitness 32
`define TB_ITERATIONS 100
