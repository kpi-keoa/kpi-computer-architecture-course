// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 64-Bit Version 13.0 (Build Build 232 06/12/2013)
// Created on Sat Sep 14 18:19:48 2019

`timescale 1 ps / 1ps

module lab2_tb;
	reg i_clk_sig;
	reg i_arst_sig;
	reg [31:0] data_sig;
	reg [4:0] adr1_sig;
	reg [4:0] adr2_sig;
	reg we_sig;
	reg [4:0] sel_sig;
	wire [31:0] Doutput1_sig;
	wire [31:0] Dout_sig;	

Block2 Block2_inst(
	.i_clk(i_clk_sig) ,	// input  i_clk_sig
	.i_arst(i_arst_sig) ,	// input  i_arst_sig
	.data(data_sig) ,	// input [31:0] data_sig
	.adr1(adr1_sig) ,	// input [4:0] adr1_sig
	.adr2(adr2_sig) ,	// input [4:0] adr2_sig
	.we(we_sig) ,	// input  we_sig
	.sel(sel_sig) ,	// input [4:0] sel_sig
	.Doutput1(Doutput1_sig) ,	// output [31:0] Doutput1_sig
	.Dout(Dout_sig) 	// output [31:0] Dout_sig
);

initial begin
	i_clk_sig =1'd1;
	forever #1 i_clk_sig = ~i_clk_sig;
end

initial begin
	i_arst_sig = 1'b1;
	we_sig = 1'b1;
	 
	#2 i_arst_sig = 1'b0;
	#2 i_arst_sig = 1'b1;
	
end



initial begin
	data_sig = 32'h0;
	forever #5 data_sig = data_sig + 1'h1;

end 

initial begin 
	adr1_sig = 5'b00000;
	adr2_sig = 5'b00000;
	
	forever #20 adr1_sig = adr1_sig + 5'h1;
	
end 

initial begin 
	sel_sig = 5'b00000;
	
	 forever #20 sel_sig = sel_sig + 5'h1;

end

initial begin
	#620 $stop();

end

endmodule
	
