// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 64-Bit Version 13.0 (Build Build 232 06/12/2013)
// Created on Mon Sep 23 21:51:54 2019
`timescale 1ns/1ps

module laba2_tb;
	reg i_we_sig;	
	reg i_clk_sig;	
	reg i_arst_sig;
	reg [4:0] WAddr_sig;	
	reg [31:0] i_d_sig; 
	reg [4:0] ReadAddrA_sig;
	reg [4:0] ReadAddrB_sig;
	wire [31:0] o_A_sig;
	wire [31:0] o_B_sig;

laba2 laba2_inst
(
	.i_we(i_we_sig) ,	// input  i_we_sig
	.i_clk(i_clk_sig) ,	// input  i_clk_sig
	.i_arst(i_arst_sig) ,	// input  i_arst_sig
	.WAddr(WAddr_sig) ,	// input [4:0] WAddr_sig
	.i_d(i_d_sig) ,	// input [31:0] i_d_sig
	.ReadAddrA(ReadAddrA_sig) ,	// input [4:0] ReadAddrA_sig
	.ReadAddrB(ReadAddrB_sig) ,	// input [4:0] ReadAddrB_sig
	.o_A(o_A_sig) ,	// output [31:0] o_A_sig
	.o_B(o_B_sig) 	// output [31:0] o_B_sig
);
	initial begin
		 i_clk_sig = 1'b0;
		 forever #10 i_clk_sig=~i_clk_sig;
		end
	
	initial begin 
		i_arst_sig=1'b1;
		#5 i_arst_sig=1'b0;
		#5 i_arst_sig=1'b1;
		end

	initial begin 
		i_d_sig=32'h11111111;		
		i_we_sig=1'b0;
		WAddr_sig = 5'b00001;
		ReadAddrA_sig=5'b00001;
		ReadAddrB_sig=5'b00000;
		#25 i_we_sig=1'b1;
		#20 i_we_sig=1'b0;
		i_d_sig=32'h33333333;
		WAddr_sig = 5'b00011;
		ReadAddrA_sig=5'b00001;
		ReadAddrB_sig=5'b00011;
		#20 i_we_sig=1'b1;
		#15 i_we_sig=1'b0;
		i_d_sig=32'h88888888;
		WAddr_sig = 5'b01000;
		ReadAddrA_sig=5'b01000;
		ReadAddrB_sig=5'b00001;
		#25 i_we_sig=1'b1;
		#15 i_we_sig=1'b0;
				
	end

	initial begin 
			#130 $stop();
	end

	endmodule
